
module negB(b, s);
    input [7:0]b;
    output [7:0]s;

    assign s = -b;

endmodule