
module negA(a, s);
    input [7:0]a;
    output [7:0]s;

    assign s = -a;

endmodule